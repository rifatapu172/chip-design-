module stimulus;
  reg I0,I1,I2,I3,S1,S0;
  wire OUT;
  mux m1(OUT,I0,I1,I2,I3,S1,S0);
  initial
  $monitor($time, "OUT=%b,S1%b=,S0=%b",OUT,S1,S0);

  initial
  begin
      I0=1'b1; I1=1'b0; I2=1'b1; I3=1'b0;
         S1=1'b0; S0=1'b0;
      #5 S1=1'b0;S0=1'b1;
      #5 S1=1'b1;S0=1'b0;
      #5 S1=1'b1;S0=1'b1;
      #5 $stop;
    end
    endmodule
